//
// Verilog Module ECC_ENC_DEC_lib.APB_SLAVE
//
// Created:
//          by - yossi.UNKNOWN (LAPTOP-LDM4S6RE)
//          at - 12:22:15 11/23/2021
//
// using Mentor Graphics HDL Designer(TM) 2018.2 (Build 19)
//

`resetall
`timescale 1ns/10ps
module APB_SLAVE ;


// ### Please start your Verilog code here ### 

endmodule
